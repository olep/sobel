-- filename: sobel.vhd
-- date: 26.08.2016

----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use sobel_package.all;
----------------------------------------------------------------------------
entity sobel is
	port (
		clk : in std_logic;
		rst : in std_logic; 
		
		
	);
end entity;
----------------------------------------------------------------------------
architecture rtl of sobel is
begin

end architecture;
----------------------------------------------------------------------------

