----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use image_proc_package.all;
----------------------------------------------------------------------------
entity image_proc_controller is
	port (
		clk : in std_logic;
		rst : in std_logic; 
		
		
	);
end entity;
----------------------------------------------------------------------------
architecture rtl of sobel_controller is
begin

end architecture;
----------------------------------------------------------------------------

